// Submit this file with other files you created.
// Do not touch port declarations of the module 'cpu'.

// Guidelines
// 1. It is highly recommened to `define opcodes and something useful.
// 2. You can modify the module.
// (e.g., port declarations, remove modules, define new modules, ...)
// 3. You might need to describe combinational logics to drive them into the module (e.g., mux, and, or, ...)
// 4. `include files if required

module cpu(input reset,                     // positive reset signal
           input clk,                       // clock signal
           output is_halted,                // Whehther to finish simulation
           output [31:0] print_reg [0:31]); // TO PRINT REGISTER VALUES IN TESTBENCH (YOU SHOULD NOT USE THIS)
    /***** declarations *****/
    // 1. pc
    
    wire [31:0] nextpcValue;
    wire [31:0] pcValue; //use this

    // 2. instruction_memory

    wire [31:0] instOutput;
    // 3. register_file
    wire [4:0] rs1, rs2, rd;
    wire [31:0] rd_din;
    wire write_enable;
    wire [31:0] rs1_dout, rs2_dout;

    // 4. control_unit

    // 5. imm gen
    wire [31:0] immgenOutput;
    // 6. alu_control_unit

    // 7. alu
    wire [2:0] alu_op;
    wire [31:0] alu_in_1, alu_in_2, alu_result;
    wire alu_bcond;

    //8. etc
    
    wire [31:0] adder1Output;
    wire [31:0] adder2Output;
    wire [31:0] mux1Output;
    wire [31:0] mux2Output;
    wire [31:0] mux3Output;
    wire [31:0] mux4Output;
    wire [31:0] mux5Output;


  /***** Wire declarations *****/
  /***** Register declarations *****/

  // ---------- Update program counter ----------
  // PC must be updated on the rising edge (positive edge) of the clock.
  pc pc(
    .reset(),       // input (Use reset to initialize PC. Initial value must be 0)
    .clk(),         // input
    .next_pc(),     // input
    .current_pc(pcValue)   // output
  );

  
  // ---------- Instruction Memory ----------
  instruction_memory imem(
    .reset(reset),   // input
    .clk(clk),     // input
    .addr(pcValue),    // input
    .dout(instOutput)     // output
  );

  // ---------- Register File ----------
  register_file reg_file (
    .reset(reset),        // input
    .clk(clk),          // input
    .rs1(rs1),          // input
    .rs2(rs1),          // input
    .rd(rd),           // input
    .rd_din(rd_din),       // input
    .write_enable(write_enable), // input
    .rs1_dout(rs1_dout),     // output
    .rs2_dout(rs2_dout),     // output
    .print_reg(print_reg)  //DO NOT TOUCH THIS
  );


  // ---------- Control Unit ----------
  control_unit ctrl_unit (
    .part_of_inst(),  // input
    .is_jal(),        // output
    .is_jalr(),       // output
    .branch(),        // output
    .mem_read(),      // output
    .mem_to_reg(),    // output
    .mem_write(),     // output
    .alu_src(),       // output
    .write_enable(),  // output
    .pc_to_reg(),     // output
    .is_ecall()       // output (ecall inst)
  );

  // ---------- Immediate Generator ----------
  immediate_generator imm_gen(
    .part_of_inst(instOutput),  // input
    .imm_gen_out(immgenOutput)    // output
  );

  // ---------- ALU Control Unit ----------
  alu_control_unit alu_ctrl_unit (
    .part_of_inst(),  // input
    .alu_op()         // output
  );

  // ---------- ALU ----------
  alu alu (
    .alu_op(alu_op),      // input
    .alu_in_1(alu_in_1),    // input  
    .alu_in_2(alu_in_2),    // input
    .alu_result(alu_result),  // output
    .alu_bcond(alu_bcond)    // output
  );

  // ---------- Data Memory ----------
  data_memory dmem(
    .reset(),      // input
    .clk(),        // input
    .addr(),       // input
    .din(),        // input
    .mem_read(),   // input
    .mem_write(),  // input
    .dout()        // output
  );

  adder adder1(
    .x1(pcValue),
    .x2(32'b100),
    .y(adder1Output)
  );

  adder adder2(
    .x1(pcValue),
    .x2(immgenOutput),
    .y(adder2Output)
  );
  2x1mux 2x1mux1(
    .x0(adder1Output),
    .x1(adder2Output),
    .sel(pcsrc1),
    .y(mux1Output)
  );
  2x1mux 2x1mux2(
    .x0(),
    .x1(),
    .sel(),
    .y()
  );
  2x1mux 2x1mux3(
    .x0(),
    .x1(immgenOutput),
    .sel(),
    .y()
  );
  2x1mux 2x1mux4(
    .x0(),
    .x1(),
    .sel(),
    .y()
  );
  2x1mux 2x1mux5(
    .x0(),
    .x1(),
    .sel(),
    .y()
  );
endmodule
